module main

import net.websocket

fn main() {
	
}

